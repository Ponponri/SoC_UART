`timescale  1ns/1ps


module split_tb;


reg [17*8:0] dict [0:62];

file = fopen('inst_matmul.dat', 'wb');
for i


endmodule